--TODO: CPU , Y MEMORIA 

--BLOQUE MEMORIA

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Practica_CIP is
  port
  (
    --entradas y salidas 

  );
end entity Practica_CIP;

architecture arch_Practica_CIP of Practica_CIP is
  
  
  -- SIGNALS --------------------------------------

begin
  

end;
-------------------------------------------   