-- 3 registros para operaciones. 2 de valores y 1 de reultados 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity alu is
  port
  (
    --entradas y salidas 
    
  );
end entity alu;

architecture arch_alu of alu is
  
    -- SIGNALS --------------------------------------
  
  
  
    -- Componentes -----------------------------------
  
  
  
  begin
    -- Instanciacion de componentes  ----------------------------
  
    
  
    -- PROCESOS --------------------------------------------------
  
  end;
  