-- Códgio de memoria definido en el enunciado de la práctica.