

--Maquina de estados

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity control_unit is
  port
  (
    --entradas y salidas 

  );
end entity control_unit;

architecture arch_control_unit of control_unit is
  
  
  -- SIGNALS --------------------------------------

begin
  

end;
-------------------------------------------   